module memory_to_reg ( 
    input [31:0] i_memory_data,
    input [31:0] i_alu_result,
    input [5:0] i_opcode,
    output reg [31:0] o_wb_data
)


endmodule
