module alu_ctrl (
    input [5:0] i_opcode,
    output reg [2:0] o_alu_ctrl
);