module sign_extend (
    input i_adress,
    input i_se_ctrl, //control signal for sign extend
    output o_extended_adress
);