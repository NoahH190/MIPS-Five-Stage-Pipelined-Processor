module shift_mux ( //shifts 5 bits 
    input i_sel_shift,
    input [4:0] i_shamt, //figure out where im pulling shampt from
    input [31:0] i_src1,
    output reg [4:0] o_shamt
);

endmodule
