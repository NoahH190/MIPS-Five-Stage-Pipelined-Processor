module shift_mux ( //shifts 5 bits 
    input i_sel_shift,
    input i_shampt, //figure out where im pulling shampt from
    input tbd,
    output reg [4:0] o_shamt
);

endmodule
