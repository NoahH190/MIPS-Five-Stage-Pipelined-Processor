module pcjump_mux (
    input i_clk,
    input i_reset,
    input i_pc_jmp_sel,
);