module and_gate (
    input i_opcode, 
    input i_zero,
    output reg o_and
)



endmodule