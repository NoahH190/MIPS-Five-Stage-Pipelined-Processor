module sign_extend (
    input [15:0] i_address,
    input i_se_ctrl, //control signal for sign extend
    output reg [21:0] o_extended_adress
);



endmodule
 
