module pcbranch_mux (
    input i_clk,
    input i_reset,
    input i_pc_br_sel,
);