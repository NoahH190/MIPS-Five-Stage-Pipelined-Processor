module alu_mux (
    input [5:0] i_sel_alu,
    input [31:0] i_sign_extend,
    input [31:0] i_src2,
    output reg [31:0] o_alu_mux
);

endmodule

