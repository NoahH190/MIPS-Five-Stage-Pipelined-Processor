module pcbranch_mux (
    input i_clk,
    input i_reset,
    input i_pc_br_sel,
    input [31:0] i_branch_adress_0,
    input [31:0] i_add_next, 
    output [31:0] o_branch_address_1
);