module sign_extend (
    input [15:0] i_address,
    input [5:0] i_se_ctrl, //control signal for sign extend
    output reg [31:0] o_sign_extend
);

endmodule
 
