module add_brn (
    input [31:0] i_address,
    input [31:0] i_add_next,
    input i_se_crtl,
    output reg [31:0] o_br_address
);


endmodule
