module data_memory(
    input i_clk,
    input i_read, //read signal
    input i_write, //write signal 
    input [31:0] tbd,   //should be output of ALU unit
    input [31:0] tbd,   //should be source 2 but have to confirm
    output reg [31:0] tbd
);

//this is most likely gonna be implemented on ddr3 ram 

endmodule 